// +FHDR----------------------------------------------------------------------------
// Project Name  : RISC-V
// Author        : shaoxuan
// Email         : caisegou@foxmail.com
// Created On    : 2023/09/18 22:34
// Last Modified : 2023/09/18 22:34
// File Name     : regfile.v
// Description   :
//         
// 
// ---------------------------------------------------------------------------------
// Modification History:
// Date         By              Version                 Change Description
// ---------------------------------------------------------------------------------
// 2023/09/18   shaoxuan        1.0                     Original
// -FHDR----------------------------------------------------------------------------
module REGFILE
(
    input       sclk_i,
    input       srst_i,

);




endmodule

